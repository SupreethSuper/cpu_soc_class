`include "regfile_defines.vh"
localparam REG_BASE_ADDR = `REG_BASE_ADDR_DEF;
localparam REG_NUM_WORDS = `REG_NUM_WORDS_DEF;
localparam REG_NUM_BITS  = `REG_NUM_BITS_DEF;

