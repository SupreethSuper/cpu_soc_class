`include "memory_defines.vh"
localparam MEM_BASE_ADDR = `MEM_BASE_ADDR_DEF;
localparam MEM_NUM_WORDS = `MEM_NUM_WORDS_DEF;
localparam MEM_NUM_BITS  = `MEM_NUM_BITS_DEF;
