`ifndef REG_DEFINES
`define REG_DEFINES

// Register-file default base address (32-bit), number of words, and bits per word
`define REG_BASE_ADDR_DEF 32'h00002000
`define REG_NUM_WORDS_DEF 32
`define REG_NUM_BITS_DEF 32

`endif // REG_DEFINES
