`ifndef MEM_DEFINES
`define MEM_DEFINES

// Memory default base address (32-bit), number of words, and bits per word
`define MEM_BASE_ADDR_DEF 32'h00001000
`define MEM_NUM_WORDS_DEF 1024
`define MEM_NUM_BITS_DEF 32

`endif // MEM_DEFINES
