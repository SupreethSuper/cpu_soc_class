`include "memory_defines.vh"

// These are localparams intended to be included inside a module or top-level
// and used for instantiation parameters / checks.
localparam MEM_BASE_ADDR  = `MEM_BASE_ADDR_DEF;
localparam MEM_NUM_WORDS  = `MEM_NUM_WORDS_DEF;
localparam MEM_NUM_BITS   = `MEM_NUM_BITS_DEF;
