localparam ADD   = 12'h020;   // done
localparam ADDI  = 12'h200;   // done
localparam ADDIU = 12'h240;   // done
localparam ADDU  = 12'h021;   // done
localparam AND   = 12'h024;   // done
localparam ANDI  = 12'h300;   // done
localparam BEQ   = 12'h100;   // done
localparam BNE   = 12'h140;   // done
localparam LW    = 12'h8C0;   // done
localparam NOR   = 12'h027;   // done
localparam OR    = 12'h025;   // done
localparam ORI   = 12'h340;   // done
localparam SLL   = 12'h000;   // done
localparam SRL   = 12'h002;   // done
localparam SW    = 12'hAC0;   // done
localparam SUB   = 12'h022;   // done
localparam SUBU  = 12'h023;   // done
localparam SRA   = 12'h003;   // done
localparam J     = 12'h080;   
localparam JAL   = 12'h0C0;   
localparam JR    = 12'h008;
localparam LBU   = 12'h900;   
localparam LHU   = 12'h940;   
localparam LL    = 12'hC00;   
localparam LUI   = 12'h3C0;   
localparam SB    = 12'hA00;   
localparam SC    = 12'hE00;   
localparam SH    = 12'hA40;   
localparam SLT   = 12'h02A;
localparam SLTI  = 12'h280;
localparam SLTIU = 12'h2C0;
localparam SLTU  = 12'h02B;
localparam HALT  = 12'hFC0;
