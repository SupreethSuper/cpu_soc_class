`include "regfile_defines.vh"

// These are localparams intended to be included inside a module or top-level
// and used for instantiation parameters / checks.
localparam REG_BASE_ADDR  = `REG_BASE_ADDR_DEF;
localparam REG_NUM_WORDS  = `REG_NUM_WORDS_DEF;
localparam REG_NUM_BITS   = `REG_NUM_BITS_DEF;
