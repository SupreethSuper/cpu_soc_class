`ifndef REG_DEFINES
`define REG_DEFINES

`define REG_BASE_ADDR_DEF 32'h2000
`define REG_NUM_WORDS_DEF 32
`define REG_NUM_BITS_DEF  32

`endif 

